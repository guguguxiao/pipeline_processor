module Alu(
    input [`ALU_OP_LENGTH] aluOpE,
    input [`WORD_WIDTH]    SrcA,
    input [`WORD_WIDTH]    SrcB,
    output [`WORD_WIDTH]   aluOutE
    );



endmodule