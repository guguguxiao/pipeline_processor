`timescale 1ns / 1ps
`include "defines.vh"

module control_unit(
         input wire                         rst,
         input wire[5:0]                    opcode, // Instruction opcode
         input wire[5:0]                    func,   // R-Type instruction function
         input wire                         isRsRtEq,

         output wire                        Regfile_weD,
         output wire                        DataMem_weD,
         output wire[`EXT_OP_LENGTH]        extOpD,
         output wire[`NPC_OP_LENGTH]        npcOp,
         output wire[`ALU_OP_LENGTH]        aluOpD,
         output wire                        aluSrc2_muxD,
         output wire[`REG_SRC_LENGTH]       regSrc_muxD,
         output wire[`REG_DST_LENGTH]       regDst_muxD,
         output wire                        memToRegD // 是否为从内存加载到寄存器中的指令
       );


// TODO
endmodule